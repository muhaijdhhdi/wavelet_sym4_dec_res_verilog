`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module: fir_coeff_rom
// Description: 优化版FIR滤波器系数ROM (Q3.18格式，21位)
//              179阶对称滤波器，只存储前90个系数 (h[0]~h[89])
//
// 系数格式：Q3.18（21位有符号）
//   3位整数（含符号）+ 18位小数 = 21位
//
// 系数来源：matlab_alg_sim/test/fir_coff_binary.txt
//
// 输出格式：展平为1890位向量 (90个系数 × 21位)
//////////////////////////////////////////////////////////////////////////////////

module fir_coeff_rom #(
    parameter COEFF_WIDTH = 21,
    parameter NUM_COEFFS = 90
)(
    output wire [NUM_COEFFS*COEFF_WIDTH-1:0] coeffs  // 1890位展平向量
);

    // Q3.18格式系数（直接从fir_coff_binary.txt读取，21位二进制）
    
    // h[0] ~ h[9]
    assign coeffs[21*0  +: 21] = 21'b000000000011001101010;  // h[0]
    assign coeffs[21*1  +: 21] = 21'b000000000001010000000;  // h[1]
    assign coeffs[21*2  +: 21] = 21'b000000000001011011100;  // h[2]
    assign coeffs[21*3  +: 21] = 21'b000000000001100100111;  // h[3]
    assign coeffs[21*4  +: 21] = 21'b000000000001101011100;  // h[4]
    assign coeffs[21*5  +: 21] = 21'b000000000001101110100;  // h[5]
    assign coeffs[21*6  +: 21] = 21'b000000000001101101101;  // h[6]
    assign coeffs[21*7  +: 21] = 21'b000000000001101000100;  // h[7]
    assign coeffs[21*8  +: 21] = 21'b000000000001011110111;  // h[8]
    assign coeffs[21*9  +: 21] = 21'b000000000001010001001;  // h[9]
    
    // h[10] ~ h[19]
    assign coeffs[21*10 +: 21] = 21'b000000000000111111101;  // h[10]
    assign coeffs[21*11 +: 21] = 21'b000000000000101011000;  // h[11]
    assign coeffs[21*12 +: 21] = 21'b000000000000010100000;  // h[12]
    assign coeffs[21*13 +: 21] = 21'b111111111111111011110;  // h[13]
    assign coeffs[21*14 +: 21] = 21'b111111111111100011011;  // h[14]
    assign coeffs[21*15 +: 21] = 21'b111111111111001100001;  // h[15]
    assign coeffs[21*16 +: 21] = 21'b111111111110110111100;  // h[16]
    assign coeffs[21*17 +: 21] = 21'b111111111110100110101;  // h[17]
    assign coeffs[21*18 +: 21] = 21'b111111111110011010011;  // h[18]
    assign coeffs[21*19 +: 21] = 21'b111111111110010011111;  // h[19]
    
    // h[20] ~ h[29]
    assign coeffs[21*20 +: 21] = 21'b111111111110010011011;  // h[20]
    assign coeffs[21*21 +: 21] = 21'b111111111110011001011;  // h[21]
    assign coeffs[21*22 +: 21] = 21'b111111111110100101110;  // h[22]
    assign coeffs[21*23 +: 21] = 21'b111111111110111000000;  // h[23]
    assign coeffs[21*24 +: 21] = 21'b111111111111001111000;  // h[24]
    assign coeffs[21*25 +: 21] = 21'b111111111111101001110;  // h[25]
    assign coeffs[21*26 +: 21] = 21'b000000000000000110100;  // h[26]
    assign coeffs[21*27 +: 21] = 21'b000000000000100100010;  // h[27]
    assign coeffs[21*28 +: 21] = 21'b000000000001000000011;  // h[28]
    assign coeffs[21*29 +: 21] = 21'b000000000001011001011;  // h[29]
    
    // h[30] ~ h[39]
    assign coeffs[21*30 +: 21] = 21'b000000000001101101110;  // h[30]
    assign coeffs[21*31 +: 21] = 21'b000000000001111011011;  // h[31]
    assign coeffs[21*32 +: 21] = 21'b000000000010000001110;  // h[32]
    assign coeffs[21*33 +: 21] = 21'b000000000001111111101;  // h[33]
    assign coeffs[21*34 +: 21] = 21'b000000000001110100110;  // h[34]
    assign coeffs[21*35 +: 21] = 21'b000000000001100001100;  // h[35]
    assign coeffs[21*36 +: 21] = 21'b000000000001000110011;  // h[36]
    assign coeffs[21*37 +: 21] = 21'b000000000000100100110;  // h[37]
    assign coeffs[21*38 +: 21] = 21'b111111111111111110100;  // h[38]
    assign coeffs[21*39 +: 21] = 21'b111111111111010101100;  // h[39]
    
    // h[40] ~ h[49]
    assign coeffs[21*40 +: 21] = 21'b111111111110101100010;  // h[40]
    assign coeffs[21*41 +: 21] = 21'b111111111110000101011;  // h[41]
    assign coeffs[21*42 +: 21] = 21'b111111111101100011011;  // h[42]
    assign coeffs[21*43 +: 21] = 21'b111111111101001000110;  // h[43]
    assign coeffs[21*44 +: 21] = 21'b111111111100110111100;  // h[44]
    assign coeffs[21*45 +: 21] = 21'b111111111100110001100;  // h[45]
    assign coeffs[21*46 +: 21] = 21'b111111111100110111101;  // h[46]
    assign coeffs[21*47 +: 21] = 21'b111111111101001010011;  // h[47]
    assign coeffs[21*48 +: 21] = 21'b111111111101101001010;  // h[48]
    assign coeffs[21*49 +: 21] = 21'b111111111110010011010;  // h[49]
    
    // h[50] ~ h[59]
    assign coeffs[21*50 +: 21] = 21'b111111111111000110011;  // h[50]
    assign coeffs[21*51 +: 21] = 21'b000000000000000000010;  // h[51]
    assign coeffs[21*52 +: 21] = 21'b000000000000111101011;  // h[52]
    assign coeffs[21*53 +: 21] = 21'b000000000001111010100;  // h[53]
    assign coeffs[21*54 +: 21] = 21'b000000000010110011101;  // h[54]
    assign coeffs[21*55 +: 21] = 21'b000000000011100101000;  // h[55]
    assign coeffs[21*56 +: 21] = 21'b000000000100001010111;  // h[56]
    assign coeffs[21*57 +: 21] = 21'b000000000100100010011;  // h[57]
    assign coeffs[21*58 +: 21] = 21'b000000000100101000100;  // h[58]
    assign coeffs[21*59 +: 21] = 21'b000000000100011011110;  // h[59]
    
    // h[60] ~ h[69]
    assign coeffs[21*60 +: 21] = 21'b000000000011111011100;  // h[60]
    assign coeffs[21*61 +: 21] = 21'b000000000011001000001;  // h[61]
    assign coeffs[21*62 +: 21] = 21'b000000000010000011000;  // h[62]
    assign coeffs[21*63 +: 21] = 21'b000000000000101111001;  // h[63]
    assign coeffs[21*64 +: 21] = 21'b111111111111010000001;  // h[64]
    assign coeffs[21*65 +: 21] = 21'b111111111101101010111;  // h[65]
    assign coeffs[21*66 +: 21] = 21'b111111111100000101001;  // h[66]
    assign coeffs[21*67 +: 21] = 21'b111111111010100100110;  // h[67]
    assign coeffs[21*68 +: 21] = 21'b111111111001010000011;  // h[68]
    assign coeffs[21*69 +: 21] = 21'b111111111000001110011;  // h[69]
    
    // h[70] ~ h[79]
    assign coeffs[21*70 +: 21] = 21'b111111110111100100101;  // h[70]
    assign coeffs[21*71 +: 21] = 21'b111111110111011000100;  // h[71]
    assign coeffs[21*72 +: 21] = 21'b111111110111101110010;  // h[72]
    assign coeffs[21*73 +: 21] = 21'b111111111000101001000;  // h[73]
    assign coeffs[21*74 +: 21] = 21'b111111111010001010011;  // h[74]
    assign coeffs[21*75 +: 21] = 21'b111111111100010010011;  // h[75]
    assign coeffs[21*76 +: 21] = 21'b111111111110111111011;  // h[76]
    assign coeffs[21*77 +: 21] = 21'b000000000010001101111;  // h[77]
    assign coeffs[21*78 +: 21] = 21'b000000000101111001000;  // h[78]
    assign coeffs[21*79 +: 21] = 21'b000000001001111010001;  // h[79]
    
    // h[80] ~ h[89]
    assign coeffs[21*80 +: 21] = 21'b000000001110001001111;  // h[80]
    assign coeffs[21*81 +: 21] = 21'b000000010010011111011;  // h[81]
    assign coeffs[21*82 +: 21] = 21'b000000010110110001101;  // h[82]
    assign coeffs[21*83 +: 21] = 21'b000000011010110111001;  // h[83]
    assign coeffs[21*84 +: 21] = 21'b000000011110100111000;  // h[84]
    assign coeffs[21*85 +: 21] = 21'b000000100001111000011;  // h[85]
    assign coeffs[21*86 +: 21] = 21'b000000100100100011111;  // h[86]
    assign coeffs[21*87 +: 21] = 21'b000000100110100011001;  // h[87]
    assign coeffs[21*88 +: 21] = 21'b000000100111110001011;  // h[88]
    assign coeffs[21*89 +: 21] = 21'b000000101000001011110;  // h[89] (中心系数)

endmodule
